A15 - LED_1
A14 - LED_2
A13 - LED_3
A12 - LED_4
E17 - LED_5


