-- pass one token between two boards
